module Testing(
 input       Clk,       // N14 = 50 MHz
 output [0:0]LVDS_TX_P, // LVDS: V17-W17

 input  [4:1]Button,    // AB5  V5 R1 M1
 output [8:1]LED        // AA5 AB4 T6 V4 T1 R2 N1 M2
);
//------------------------------------------------------------------------------

assign LED       = {Button, Button};
assign LVDS_TX_P = Clk;
//------------------------------------------------------------------------------

endmodule
//------------------------------------------------------------------------------
 