module Testing(
 input  Clk,
 output [0:0]LVDS_TX_P,
 input  [4:1]Button,
 output [8:1]LED
);
//------------------------------------------------------------------------------

assign LED = {2{Button}};
assign LVDS_TX_P = Clk;
assign Testing = 16'hABCD;
//------------------------------------------------------------------------------

endmodule
//------------------------------------------------------------------------------

